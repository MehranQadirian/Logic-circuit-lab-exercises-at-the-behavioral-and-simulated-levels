`timescale 1ns / 1ps
module Multiplier4x3 (
    input [3:0] A,
    input [2:0] B,
    output [6:0] Y
);
    // ?????????? ????? ???? ??????? ????
    wire [3:0] partial_prod [2:0];
    wire [3:0] sum [1:0];
    wire [1:0] carry;

    // ?????? ??????????? ????
    assign partial_prod[0] = {4{B[0]}} & A;  // A * B[0]
    assign partial_prod[1] = {4{B[1]}} & A;  // A * B[1]
    assign partial_prod[2] = {4{B[2]}} & A;  // A * B[2]

    // ????????????? ? ???? ???? ??????? ????
    FullAdder4bit FA1 (
        .A({1'b0, partial_prod[0][3:1]}),
        .B(partial_prod[1]),
        .C_in(1'b0),
        .Sum(sum[0]),
        .C_out(carry[0])
    );

    FullAdder4bit FA2 (
        .A({carry[0], sum[0][3:1]}),
        .B(partial_prod[2]),
        .C_in(1'b0),
        .Sum(sum[1]),
        .C_out(carry[1])
    );

    // ????? ????? ?????
    assign Y = {carry[1], sum[1], sum[0][0], partial_prod[0][0]};
endmodule