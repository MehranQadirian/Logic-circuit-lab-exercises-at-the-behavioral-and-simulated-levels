`timescale 1ns / 1ps

module main(
    input A, B, C, D,
    output F1, F2
);
    // ????? ??????? ????
    wire T1, T2, T3, T4;

    // ?????? ??????? ???? ?? ???? ????????
    assign T1 = A & B;   // T1 = AND(A, B)
    assign T2 = B | C;   // T2 = OR(B, C)
    assign T3 = C ^ D;   // T3 = XOR(C, D)
    assign T4 = ~D;      // T4 = NOT(D)

    // ?????? ????????? ????? ?? ???? ??????? ????
    assign F1 = T1 | T3; // F1 = OR(T1, T3)
    assign F2 = T2 & T4; // F2 = AND(T2, T4)

endmodule
