
`timescale 1ns / 1ps

module FourBitAdder_TB;  // ??? ?????????
    reg [3:0] A, B;
    reg C_in;
    wire [3:0] S;
    wire C_out, V;
    
    // ???????? ?? ???? ????
    FourBitAdder uut (
        .A(A),
        .B(B),
        .C_in(C_in),
        .S(S),
        .C_out(C_out),
        .V(V)
    );
    
    initial begin
        // ??????? ?????
        A = 4'b0010; B = 4'b0001; C_in = 0;  // ??? ?: 2 + 1
        #10;
        
        A = 4'b1000; B = 4'b1000; C_in = 0;  // ??? ?: 8 + 8 (????? ???? ?????)
        #10;
        
        A = 4'b0111; B = 4'b0001; C_in = 0;  // ??? ?: 7 + 1 (????? ?????????)
        #10;
        
        A = 4'b1111; B = 4'b0000; C_in = 1;  // ??? ?: 15 + 0 + 1 (??? Carry-in)
        #10;
        
    end
endmodule